`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Description: 1λ�ӷ�������32λcla��ײ��ģ��
//              ���룺����1λ����a,b��һ����λ��λc
//              �����1λ�ӷ����s����λ��������g����λ���ݺ���p
//////////////////////////////////////////////////////////////////////////////////


module add_1 (a,b,c, g,p,s);
    input a,b,c;
    output g,p,s;
    assign s = a ^ b ^ c;
    assign g = a & b;
    assign p = a | b;
endmodule
