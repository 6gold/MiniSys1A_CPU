`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Description: 
//////////////////////////////////////////////////////////////////////////////////

module MinisysEXE(
    //input
    clk,rst,control,srca,srcb,shamt,immi,hi2regdata,lo2regdata,mfc0data,pc_in,intr,runoverflow,icmisspause,dcmisspause,dtlbRefill_exc,
    //output
    exepwreg,exepmem2reg,exepwaddreg,exepalu,exeresult,exewmdata,execontrol,overflow,                                          
    prerror,mulbusy,divbusy,keepmd,mulover,divover,exepmdcs,exepmdhidata,exepmdlodata,exemdhidata,exemdlodata,exemdcs,         //output
    /*md,*/exebranch,pctoid,exetomempc);
    
    //�����������
    /* ��ALU��ص� */
    //sub_add
    //�߼�����
    
    
    
    /* ��ALU��ص� */
    //mult_div
    
    
    
    //������ѡ��
endmodule
